--FPQ.VHD
           LIBRARY IEEE;
           USE IEEE.STD_LOGIC_1164.ALL;
           USE IEEE.STD_LOGIC_UNSIGNED.ALL;
           USE IEEE.STD_LOGIC_ARITH.ALL;
           ENTITY FPQ IS
PORT(SCLK: IN STD_LOGIC;    		--SCLK=200 Hz
	       CLK1HZ: OUT STD_LOGIC); --CLK1HZ=1 Hz
END ENTITY FPQ; 
ARCHITECTURE ART OF FPQ IS
  SIGNAL CNT100: INTEGER RANGE 0 TO 99; 
  SIGNAL CLK1: STD_LOGIC;
  BEGIN
  PROCESS(SCLK)
BEGIN
    IF SCLK'EVENT AND SCLK='1' THEN
	      IF CNT100=99 THEN     
	        CNT100<=0;
	        CLK1<=NOT CLK1;
	      ELSE 
	        CNT100<=CNT100+1;
	      END IF;
    ELSE 
CLK1<=CLK1;
    END IF;
    CLK1HZ<=CLK1;
  END PROCESS;
END ARCHITECTURE ART;
