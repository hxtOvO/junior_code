--DDPB.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY DDPB IS
  PORT(START,WCLK:IN STD_LOGIC;
	   CLK1HZ:IN STD_LOGIC;  
	   DDBZ:OUT STD_LOGIC); 
END ENTITY DDPB;
ARCHITECTURE ART OF DDPB IS
  SIGNAL T60S:STD_LOGIC;  
  SIGNAL WCLKCOU:STD_LOGIC_VECTOR(7 DOWNTO 0);  
  BEGIN
  --����60 s�����������źŽ���
  PROCESS(START, CLK1HZ) IS
    VARIABLE CNT60: STD_LOGIC_VECTOR(7 DOWNTO 0);
    BEGIN
    IF START='1' THEN
CNT60:="00000000"; T60S<='0';
    ELSIF CLK1HZ'EVENT AND CLK1HZ='1' THEN
      IF CNT60="00111100" THEN --CNT60=60
  	    T60S<='1'; CNT60:="00000000";
  	  ELSE
  	    CNT60:=CNT60+'1'; T60S<='0';
      END IF; 
    END IF; 
  END PROCESS ;
  --ÿ������ʻ����������
PROCESS(START, WCLK, T60S) IS
    BEGIN
    IF START='1' THEN
      WCLKCOU<="00000000";
    ELSIF WCLK'EVENT AND WCLK='1' THEN
      IF T60S='1' THEN 
        WCLKCOU<="00000000";
      ELSE
	        WCLKCOU<=WCLKCOU+'1';	
                                            --������㣬��λΪm
END IF; 
    END IF;
  END PROCESS ;
  --�ȴ���־�б����
  PROCESS(WCLKCOU,T60S) IS 
    BEGIN
    IF T60S'EVENT AND T60S='1' THEN 
      IF WCLKCOU<="11001000" THEN --WCLKCOU<=200 
	    DDBZ<='1';  --�ȴ�
      ELSE
DDBZ<='0';  --��ʻ
      END IF; 
    END IF;
  END PROCESS ; 
END ARCHITECTURE ART;

