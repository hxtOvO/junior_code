--DDJS.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY DDJS IS
  PORT(START, DDBZ: IN STD_LOGIC;
	       CLK1HZ: IN STD_LOGIC;
	       DDSJ: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);

XDBZ: OUT STD_LOGIC);
END ENTITY DDJS;
ARCHITECTURE ART OF DDJS IS
  SIGNAL MS,MG,FS, FG: STD_LOGIC_VECTOR(3 DOWNTO 0);
  SIGNAL XIDENG: STD_LOGIC;	
  BEGIN 
  PROCESS(START, DDBZ, CLK1HZ) IS 
    BEGIN
    IF START='1' THEN
MS<="0000";MG<="0000";
	      FS<="0000";FG<="0000";
    ELSIF CLK1HZ'EVENT AND CLK1HZ='1' THEN
      IF DDBZ='1' THEN
	        IF MG=9 THEN MG<="0000";
		      IF MS=5 THEN MS<="0000";
		        IF FG=9 THEN FG<="0000";
			      IF FS=5 THEN
                XIDENG<='1';FS<="0000";
			  ELSE
FS<=FS+'1';    	--����ʮλ����      	
			  END IF;
		    ELSE
            FG<=FG+'1';   	--������λ����
		    END IF;
	      ELSE
          MS<=MS+'1';    	--����ʮλ����
	      END IF;
	    ELSE
        MG<=MG+'1';      	--������λ����

END IF;
      END IF;
    END IF;
  END PROCESS;
  XDBZ<=XIDENG;
  DDSJ(15 DOWNTO 12)<=FS;
  DDSJ(11 DOWNTO 8)<=FG;
  DDSJ(7 DOWNTO 4)<=MS;
  DDSJ(3 DOWNTO 0)<=MG;
END ARCHITECTURE ART;
