--LCJF.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY LCJF IS
  GENERIC(SD1:INTEGER:=140;   --04:00��23:00����
 		  SD2:INTEGER:=180);  --����ʱ�ε���

PORT(LCBZ,JFBZ,START,DDBZ,SDBZ:IN STD_LOGIC;
	       LCFY:OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END ENTITY LCJF;
ARCHITECTURE ART OF LCJF IS
  SIGNAL LCFY1: STD_LOGIC_VECTOR(15 DOWNTO 0);
  BEGIN
  PROCESS(START, LCBZ, SDBZ, JFBZ)
    BEGIN
    IF START='1' THEN
LCFY1<="0000000000000000";
    ELSIF JFBZ'EVENT AND JFBZ='1' THEN
      IF DDBZ='0' THEN  		--��ʻ״̬
        IF LCBZ='0' THEN    		--2 km����
	          LCFY1<="0000000000000000";
        ELSIF LCBZ='1' THEN 		--2 km����
	          IF SDBZ='0' THEN
	            LCFY1<=LCFY1+SD1;
          ELSIF SDBZ='1' THEN
	            LCFY1<=LCFY1+SD2;
	          END IF;
END IF;
      END IF;
    END IF;
  END PROCESS;
  LCFY<=LCFY1;
END ARCHITECTURE ART;

